module userInput(Clock, Reset, 